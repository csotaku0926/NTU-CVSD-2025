// list all paths to your design files
`include "../sram_512x8/sram_512x8.v"
`include "../01_RTL/core.v"
